
module hello_world (
	clk_clk,
	reset_reset_n,
	switch_external_connection_export,
	led_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	input		switch_external_connection_export;
	output		led_external_connection_export;
endmodule
