
// This verilog file describes a synchronous n-bit counter circuit with an asynchronous, active low reset. This counter will go up until k-1, then rollover and indicate such with the rollover bit

module counter (Clock, Reset_n, Q, Rollover);
	parameter n = 4; 		// Quantity of bits for the counter, default = 4
	parameter k = 15;		// Highest value of counter, default = 15
	
	input Clock, Reset_n;
	output [n-1:0] Q;
	output Rollover;
	
	reg [n-1:0] Q;
	reg Rollover;
	
	always @(posedge Clock or negedge Reset_n)
	begin
		if(!Reset_n) begin		// Active low reset
			Q <= 1'b0;
			Rollover <= 1'b0;
		end else begin
			// Count up from Q = 0 to k-1
			if(Q < k-1)
			begin
				Q <= Q + 1'b1;
				Rollover <= 1'b0;
			end
			else
			begin
				Q <= 0;
				Rollover <= 1'b1;
			end
//			// Rollover (has to be k-2 due to non-blocking assignments):
//			if (Q == k-2)
//				Rollover <= 1'b1;
//			else
//				Rollover <= 1'b0;
		end
	end
endmodule